version https://git-lfs.github.com/spec/v1
oid sha256:92e7a20507234f95cd7d52d3a5b8cc55cc6320b51067222fc123da61f7dc015c
size 7712
