version https://git-lfs.github.com/spec/v1
oid sha256:d155d5a0fba179b92e034115643b80320f38e260c5de09a882e8ba191f925792
size 4640
