version https://git-lfs.github.com/spec/v1
oid sha256:3910a7f4a46408520b03824a7209a31f18555dd498477e18e0dfe2ed67d04a28
size 7712
