version https://git-lfs.github.com/spec/v1
oid sha256:4abbca0967bd36d53db848cc6e3d3532faa83f3c56777a9dce6afecdc3db0182
size 10272
