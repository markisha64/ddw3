version https://git-lfs.github.com/spec/v1
oid sha256:2d77fb0d87c52505b55d5f55f60607534f60748436253f1d66272c15005c46b7
size 8736
