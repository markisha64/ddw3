version https://git-lfs.github.com/spec/v1
oid sha256:241db082a6efd8b0a5920956a28556e7fe0ee3efa7819b71ab8ac26af8fb2d52
size 8736
