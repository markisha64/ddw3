version https://git-lfs.github.com/spec/v1
oid sha256:3ff72455afd7fbc014207b202988dbe2ab4f42d61865f1c236f80f47ef308b49
size 10272
