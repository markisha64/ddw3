version https://git-lfs.github.com/spec/v1
oid sha256:41c3079563b3faeeb3e535a2faedb3c0303bad2e37e7408b0649d3cd016ce3d3
size 9760
