version https://git-lfs.github.com/spec/v1
oid sha256:83c1bc27531bed21029f157b07857467aaebf3dde5e97eb0677ba84c33a6ce03
size 7712
