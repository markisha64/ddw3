version https://git-lfs.github.com/spec/v1
oid sha256:87944c593cb24a58547fdc9cc1d1723d285e60aee454e6ee9fcccc95da19a0c7
size 10784
