version https://git-lfs.github.com/spec/v1
oid sha256:d29695dfea4ed74d855d097e9d9e2fa7baf4019520386f0340ad9c816a5d1fc9
size 5664
