version https://git-lfs.github.com/spec/v1
oid sha256:dc444482ce08df5c972e8565e2fb32d907862c3cbec479df54cabf3d9c4b3e15
size 5152
