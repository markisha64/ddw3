version https://git-lfs.github.com/spec/v1
oid sha256:d3651264f2b7fc4fa5a265a5bdf43471f78892bc18f1a2fec75469b1669ec866
size 6688
