version https://git-lfs.github.com/spec/v1
oid sha256:15dbc227fa87a7f4776ee81291f6e2a4b313163cb03f0e59c2635da88d15e41b
size 7712
