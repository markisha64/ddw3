version https://git-lfs.github.com/spec/v1
oid sha256:4bb78b1a3d84570ed15f127117fba357a4c46d23765ff65cba6843f3e8c561f0
size 10272
