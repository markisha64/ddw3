version https://git-lfs.github.com/spec/v1
oid sha256:4851312fd5ce304a73802b72985fa3eced8c2609f423d069b642fe07066a8a0c
size 8224
