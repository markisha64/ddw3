version https://git-lfs.github.com/spec/v1
oid sha256:534fc5cab55f26fa7fc2e646161bf630accee9f0fef78a84a5c6b422adbc3d9e
size 9248
