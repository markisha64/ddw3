version https://git-lfs.github.com/spec/v1
oid sha256:790c48359bad3357734a39646d246abf968474da7a8044ffe8f3e85c92efc620
size 7712
