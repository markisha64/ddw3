version https://git-lfs.github.com/spec/v1
oid sha256:bb7ba34c36d1956f886c6e36b0cdd7240d50a1d3e44aa69fb19bcf57796c3940
size 18168
