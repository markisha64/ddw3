version https://git-lfs.github.com/spec/v1
oid sha256:6af0f6821b39f216d1a79158c9747d4a797f2e21926e9ab2af5ca9f2215355e2
size 5152
