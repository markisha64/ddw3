version https://git-lfs.github.com/spec/v1
oid sha256:c43c91a661b1da8183485a43bcf09b58c8656e1d252283c0fc50d09c1c6a5872
size 4640
