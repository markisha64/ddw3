version https://git-lfs.github.com/spec/v1
oid sha256:bf5a412e51c9749309749536b32fbe8c407f11f90875b62383374b92dc4705d6
size 7712
