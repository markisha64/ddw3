version https://git-lfs.github.com/spec/v1
oid sha256:efd92d97c95d96867fcc7133becdaa1300f028de51e705e8861ca2aef8ddde16
size 4640
