version https://git-lfs.github.com/spec/v1
oid sha256:1efeb1cc1aa7c45bb9a8f422fcb4e02ded4a8a98c5461ef5bbfe7b8e0f84fc02
size 7712
