version https://git-lfs.github.com/spec/v1
oid sha256:ab2e3d6cd7cb9705d4aac0d6df1a6f34200a2bac9ecf7680c0e31de1616104d9
size 7200
