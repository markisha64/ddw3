version https://git-lfs.github.com/spec/v1
oid sha256:0377f4a650f05f68c159ddc2454f34ab34b5faca5a096f06986c539fbd330a3e
size 8736
