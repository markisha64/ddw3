version https://git-lfs.github.com/spec/v1
oid sha256:9ab403a74ab69af9581ba1bb9b02c1b3c70ceeb8e7c6a2ba86c4508877413714
size 7200
