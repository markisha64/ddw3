version https://git-lfs.github.com/spec/v1
oid sha256:23974c73eeb8dd24968a62dc84f44e0034e7c645384c844e4bc3f6732cae5574
size 8736
