version https://git-lfs.github.com/spec/v1
oid sha256:fde7f3d2cee4df766d45d96a1c9c283c74a851b52f8db834ef57cf8c3cf02851
size 4128
