version https://git-lfs.github.com/spec/v1
oid sha256:81b8c65c11206548ae7c8cf892aa8de55b4d3f051a78d7cb44226f0d25ac737d
size 10272
