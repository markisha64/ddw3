version https://git-lfs.github.com/spec/v1
oid sha256:a2ebfcc737e6b4217d4a6b76c29dd7fe407dc2559f13b8bb694e90267f7cfee0
size 5152
