version https://git-lfs.github.com/spec/v1
oid sha256:490946c8f58a637b8ef528c29db2bcf5236581cfe80a5ace57b66d44c5cf5fab
size 8736
