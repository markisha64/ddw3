version https://git-lfs.github.com/spec/v1
oid sha256:0cc3a435e7a3ec38b2f14b6f6717302cc986bc63113f495872821292471edba5
size 4640
