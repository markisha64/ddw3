version https://git-lfs.github.com/spec/v1
oid sha256:6831a110fa68002dfcb45aed63920bce60e7968a9785b8bc1b8ba5e93a04deff
size 5152
