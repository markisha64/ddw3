version https://git-lfs.github.com/spec/v1
oid sha256:8e4b58755a8a099b12ce4078505778cd5104479e918c2fcf48a5450c3e90403a
size 4640
