version https://git-lfs.github.com/spec/v1
oid sha256:5e55860b22141b69b337ef9b8fe20d4a08940fc58b6575baab53cd3896d39d93
size 7712
